// 按键模块
module Buttons(
    
);

endmodule