// 7段数码管驱动模块
module Seg7(
    
);

endmodule